module Q_EXPLOIT (
	input logic clk,
	input logic rst,
	input logic [31:0] final_Q [37][4],
	input logic [5:0] blocked [16],
	input logic [5:0] target_state,
	input logic [5:0] start_state,
	input logic move_complete,
	input logic [5:0] maze_state,
	output logic [5:0] next_state,
	output logic timer_start);
//	output logic target_reached);
	
//	wire [5:0] blocked[16];
//	wire [31:0] final_Q [37][4];
//	wire [5:0] maze_state ;
	wire logic [31:0] max_Q;
	wire logic [3:0] action;
//	wire [31:0] reward;
	wire logic done;
	
	ACTION_EXPLOIT ACTION_EXPLOIT(
	.old_Q(final_Q), .maze_state(maze_state), .clk(clk), .rst(rst), .max_Q(max_Q), .action(action), .move_complete(move_complete), .done(done));
					
	Q_TRIAL_EXPLOIT Q_TRIAL_EXPLOIT(
	.old_Q(final_Q), .action(action), .clk(clk), .rst(rst), .maze_state(maze_state), .blocked(blocked), .next_state(next_state), .start_state(start_state), .target_state(target_state), .move_complete(move_complete), .timer_start(timer_start), .done(done));
 //.target_reached(target_reached),
	endmodule
	