module KEY_INPUT(
	input logic KEY0,
	input logic KEY3,
	input logic SW1,
	input logic SW2,
	input logic SW3,
	input logic SW4,
	output logic [7:0]angle1,
	output logic [7:0]angle2,
	output logic [7:0]angle3,
	output logic [7:0]angle4,
	output logic [11:0]angle_out);
	
	logic [3:0] switches;
	logic [3:0] out1_1, out1_2, out1_3;
	//logic [3:0] angleswitch;
	assign switches = {SW1,SW2,SW3,SW4};
	
	
	always@(posedge KEY0 or posedge KEY3)
	begin
		if (switches == 4'b1000) //1
			begin
				if (KEY0 == 1)
					angle1 = angle1+1;
				else
					angle1 = angle1-1;
				case(angle1)
					>= 100:out1_3 = 1;
					<= 100:out1_3 = 0;	
					>= 90:out1_3 = 1;	
				endcase
			end
			else if (switches == 4'b0100) //2
			begin
				if (KEY0 == 1)
					angle2 = angle2+1;
				else
					angle2 = angle2-1;
			end
			else if (switches == 4'b0010) //3
			begin
				if (KEY0 == 1)
					angle3 = angle3+1;
				else
					angle3 = angle3-1;
			end
			else if (switches == 4'b0001) //4
			begin
				if (KEY0 == 1)
					angle4 = angle4+1;
				else
					angle4 = angle4-1;
			end
	end
	
endmodule
