module Q_TRIAL_EXPLOIT(
	output logic [5:0] next_state,
	output logic timer_start,
//	output logic target_reached,
	input logic clk,
	input logic rst,
	input logic [31:0] old_Q [37][4],
	input logic [3:0] action,
	input logic [5:0] maze_state,
	input logic [5:0] blocked [16],
	input logic [5:0] target_state,
	input logic [5:0] start_state,
	input logic move_complete,
	input logic done);
	
	
	logic done_clk;
	always_ff @(clk)
	begin
		if (done == 1)
			done_clk = clk;
		else 
			done_clk = 0;
		end
		
	always@(posedge done_clk)
	begin
			if (rst == 0)
				timer_start <= 1;
			if (move_complete == 0)
				timer_start <= 1;
			else
			begin
				timer_start <= 0;
				case(action)
				default: next_state <= maze_state;
				0: begin 
						if ((maze_state + 6 <= 36) && (maze_state + 6 != blocked[0] || maze_state + 6 != blocked[1] || maze_state + 6 != blocked[2] || maze_state + 6 != blocked[3] || maze_state + 6 != blocked[4] || maze_state + 6 != blocked[5] || maze_state + 6 != blocked[6] || maze_state + 6 != blocked[7] || maze_state + 6 != blocked[8] || maze_state + 6 != blocked[9] || maze_state + 6 != blocked[10] || maze_state + 6 != blocked[11] || maze_state + 6 != blocked[12] || maze_state + 6 != blocked[13] || maze_state + 6 != blocked[14] || maze_state + 6 != blocked[15]))
							next_state <= maze_state + 6'd6;
						else
							next_state <= maze_state;
					end
				1: begin 
						if ((maze_state + 1 <= 36) && (maze_state + 1 != blocked[0] || maze_state + 1 != blocked[1] || maze_state + 1 != blocked[2] || maze_state + 1 != blocked[3] || maze_state + 1 != blocked[4] || maze_state + 1 != blocked[5] || maze_state + 1 != blocked[6] || maze_state + 1 != blocked[7] || maze_state + 1 != blocked[8] || maze_state + 1 != blocked[9] || maze_state + 1 != blocked[10] || maze_state + 1 != blocked[11] || maze_state + 1 != blocked[12] || maze_state + 1 != blocked[13] || maze_state + 1 != blocked[14] || maze_state + 1 != blocked[15] || maze_state + 1 != 7 || maze_state + 1 != 13 || maze_state + 1 != 19 || maze_state + 1 != 25 || maze_state + 1 != 31))
							next_state <= maze_state + 6'd1;
						else
							next_state <= maze_state;
					end
				2: begin 
						if ((maze_state - 6 >= 1) && (maze_state - 6 != blocked[0] || maze_state - 6 != blocked[1] || maze_state - 6 != blocked[2] || maze_state - 6 != blocked[3] || maze_state - 6 != blocked[4] || maze_state - 6 != blocked[5] || maze_state - 6 != blocked[6] || maze_state - 6 != blocked[7] || maze_state - 6 != blocked[8] || maze_state - 6 != blocked[9] || maze_state - 6 != blocked[10] || maze_state - 6 != blocked[11] || maze_state - 6 != blocked[12] || maze_state - 6 != blocked[13] || maze_state - 6 != blocked[14] || maze_state - 6 != blocked[15]))
							next_state <= maze_state - 6'd6;
						else
							next_state <= maze_state;
					end
				3: begin 
						if ((maze_state + 1 <= 36) && (maze_state - 1 != blocked[0] || maze_state - 1 != blocked[1] || maze_state - 1 != blocked[2] || maze_state - 1 != blocked[3] || maze_state - 1 != blocked[4] || maze_state - 1 != blocked[5] || maze_state - 1 != blocked[6] || maze_state - 1 != blocked[7] || maze_state - 1 != blocked[8] || maze_state - 1 != blocked[9] || maze_state - 1 != blocked[10] || maze_state - 1 != blocked[11] || maze_state - 1 != blocked[12] || maze_state - 1 != blocked[13] || maze_state - 1 != blocked[14] || maze_state - 1 != blocked[15] || maze_state - 1 != 6 || maze_state - 1 != 12 || maze_state - 1 != 18 || maze_state - 1 != 24 || maze_state - 1 != 30))
							next_state <= maze_state - 6'd1;
						else
							next_state <= maze_state;
					end
				endcase
		end
		end

//	always_ff @(negedge rst or posedge done_clk)
//		begin
//				if (rst == 0 || move_complete == 0)
//					timer_start = 1;
//				else
//				begin
//					timer_start = 0;
//					case(action)
//					default: next_state = maze_state;
//					0: begin 
//							if ((maze_state + 6 <= 36) && (maze_state + 6 != blocked[0] || maze_state + 6 != blocked[1] || maze_state + 6 != blocked[2] || maze_state + 6 != blocked[3] || maze_state + 6 != blocked[4] || maze_state + 6 != blocked[5] || maze_state + 6 != blocked[6] || maze_state + 6 != blocked[7] || maze_state + 6 != blocked[8] || maze_state + 6 != blocked[9] || maze_state + 6 != blocked[10] || maze_state + 6 != blocked[11] || maze_state + 6 != blocked[12] || maze_state + 6 != blocked[13] || maze_state + 6 != blocked[14] || maze_state + 6 != blocked[15]))
//								next_state = maze_state + 6'd6;
//							else
//								next_state = maze_state;
//						end
//					1: begin 
//							if ((maze_state + 1 <= 36) && (maze_state + 1 != blocked[0] || maze_state + 1 != blocked[1] || maze_state + 1 != blocked[2] || maze_state + 1 != blocked[3] || maze_state + 1 != blocked[4] || maze_state + 1 != blocked[5] || maze_state + 1 != blocked[6] || maze_state + 1 != blocked[7] || maze_state + 1 != blocked[8] || maze_state + 1 != blocked[9] || maze_state + 1 != blocked[10] || maze_state + 1 != blocked[11] || maze_state + 1 != blocked[12] || maze_state + 1 != blocked[13] || maze_state + 1 != blocked[14] || maze_state + 1 != blocked[15] || maze_state + 1 != 7 || maze_state + 1 != 13 || maze_state + 1 != 19 || maze_state + 1 != 25 || maze_state + 1 != 31))
//								next_state = maze_state + 6'd1;
//							else
//								next_state = maze_state;
//						end
//					2: begin 
//							if ((maze_state - 6 >= 1) && (maze_state - 6 != blocked[0] || maze_state - 6 != blocked[1] || maze_state - 6 != blocked[2] || maze_state - 6 != blocked[3] || maze_state - 6 != blocked[4] || maze_state - 6 != blocked[5] || maze_state - 6 != blocked[6] || maze_state - 6 != blocked[7] || maze_state - 6 != blocked[8] || maze_state - 6 != blocked[9] || maze_state - 6 != blocked[10] || maze_state - 6 != blocked[11] || maze_state - 6 != blocked[12] || maze_state - 6 != blocked[13] || maze_state - 6 != blocked[14] || maze_state - 6 != blocked[15]))
//								next_state = maze_state - 6'd6;
//							else
//								next_state = maze_state;
//						end
//					3: begin 
//							if ((maze_state + 1 <= 36) && (maze_state - 1 != blocked[0] || maze_state - 1 != blocked[1] || maze_state - 1 != blocked[2] || maze_state - 1 != blocked[3] || maze_state - 1 != blocked[4] || maze_state - 1 != blocked[5] || maze_state - 1 != blocked[6] || maze_state - 1 != blocked[7] || maze_state - 1 != blocked[8] || maze_state - 1 != blocked[9] || maze_state - 1 != blocked[10] || maze_state - 1 != blocked[11] || maze_state - 1 != blocked[12] || maze_state - 1 != blocked[13] || maze_state - 1 != blocked[14] || maze_state - 1 != blocked[15] || maze_state - 1 != 6 || maze_state - 1 != 12 || maze_state - 1 != 18 || maze_state - 1 != 24 || maze_state - 1 != 30))
//								next_state = maze_state - 6'd1;
//							else
//								next_state = maze_state;
//						end
//					endcase
//			end
//			end	
//	
endmodule