module ACTION_EXPLOIT (
	output logic [31:0] max_Q,
	output logic [3:0] action,
	output logic done_o,
	input logic  [31:0] old_Q [37][4],
	input logic [5:0] maze_state,
	input logic clk,
	input logic rst,
	input logic move_complete,
	input logic done,
	input logic done_t);

	logic start;
	logic [31:0] current_Q[4];
	always@(clk)
	begin
		if (done == 1)
			start = clk;
		else
			start = 0;
	end
	
	always@(posedge start)
	begin
		current_Q <= old_Q[maze_state];
		if (done_t == 1)
			done_o <= 0;
		else if (move_complete == 1 && current_Q[0] > current_Q[1] && current_Q[0] > current_Q[2] && current_Q[0] > current_Q[3])
			begin
				max_Q <= current_Q[0];
				action  <= 3'd0;
				done_o <= 1;
			end
		else if (move_complete == 1 && current_Q[1] > current_Q[0] && current_Q[1] > current_Q[2] && current_Q[1] > current_Q[3])
			begin
				max_Q <= current_Q[1];
				action  <= 3'd1;
				done_o <= 1;
			end
		else if (move_complete == 1 && current_Q[2] > current_Q[1] && current_Q[2] > current_Q[0] && current_Q[2] > current_Q[3])
			begin
				max_Q <= current_Q[2];
				action  <= 3'd2;
				done_o <=1;
			end
		else if (move_complete == 1 && current_Q[3] > current_Q[1] && current_Q[3] > current_Q[2] && current_Q[3] > current_Q[0])
			begin
				max_Q <= current_Q[3];
				action  <= 3'd3;
				done_o <=1;
			end
	end
	
	
endmodule
